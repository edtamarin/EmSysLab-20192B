/home/edian/Nextcloud/Documents/ESL/Decoder/decoder_tb_post.vhd