/home/edian/Nextcloud/Documents/ESL/Decoder/decoder.vhd