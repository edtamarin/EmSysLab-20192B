/home/edian/Nextcloud/Documents/ESL/Decoder/decoder_tb.vhd