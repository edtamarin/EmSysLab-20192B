/home/edian/Nextcloud/Documents/ESL/PWMsource/pwm.vhd